`timescale 1ns/1ps

module ID (
  input logic CLK,
  input logic RST,
  input logic [15:0] ID_IN
);
  
endmodule